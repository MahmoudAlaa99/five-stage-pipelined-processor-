LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY control_unit IS
GENERIC ( n : integer := 32);
PORT( Clk,Rst,Int: IN std_logic;
	OpCode: IN std_logic_vector(4 DOWNTO 0);
	q: OUT std_logic_vector(26 DOWNTO 0);
	RtiRet: OUT std_logic
);
END control_unit;

ARCHITECTURE a_control_unit OF control_unit IS
BEGIN

PROCESS(Clk,Rst,Int)
BEGIN
IF(Rst='1')THEN
	q <= "000000000001111100000000000";	--NOP
ELSIF(Int='1')THEN
	q <= (OTHERS=>'Z');
ELSIF rising_edge(Clk)THEN
IF (OpCode = "00000") THEN	--CLC
	q <= "000000000001111110000000000";
ELSIF (OpCode = "00001") THEN	--STC
	q <= "000000000001111111000000000";
ELSIF (OpCode = "00010") THEN	--NOP
	q <= "000000000001111100000000000";
ELSIF (OpCode = "00011") THEN	--NOT Rdst
	q <= "001100000001011100000000010";
ELSIF (OpCode = "00100") THEN	--INC Rdst
	q <= "001100000001011000000000010";
ELSIF (OpCode = "00101") THEN	--DEC Rdst
	q <= "001100000001001100000000010";
ELSIF (OpCode = "00110") THEN	--OUT Rdst
	q <= "001000000011111100000000000";
ELSIF (OpCode = "00111") THEN	--IN
	q <= "000100000001111100000000000";
ELSIF (OpCode = "01000") THEN	--SWAP
	q <= "001110000001000000000000010";	
ELSIF (OpCode = "01001") THEN	--ADD
	q <= "001100100001000100000000010";
ELSIF (OpCode = "01010") THEN	--IADD
	q <= "011100100000000100000000010";
ELSIF (OpCode = "01011") THEN	--SUB
	q <= "001100100001001000000000010";
ELSIF (OpCode = "01100") THEN	--AND
	q <= "001100100001010000000000010";
ELSIF (OpCode = "01101") THEN	--OR
	q <= "001100100001010100000000010";
ELSIF (OpCode = "01110") THEN	--SHL
	q <= "001100000001110000000000010";
ELSIF (OpCode = "01111") THEN	--SHR
	q <= "001100000001100000000000010";
ELSIF (OpCode = "10000") THEN	--PUSH
	q <= "001000000001000000010100001";
ELSIF (OpCode = "10001") THEN	--POP
	q <= "000100000001111100110010001";
ELSIF (OpCode = "10010") THEN	--LDM
	q <= "010100000001111100000000011";
ELSIF (OpCode = "10011") THEN	--LDD
	q <= "010101000001111100000010001";
ELSIF (OpCode = "10100") THEN	--STD
	q <= "011001000001000000000100001";
ELSIF (OpCode = "10101") THEN	--JZ
	q <= "001000010001111100000000010";
ELSIF (OpCode = "10110") THEN	--JN
	q <= "001000010101111100000000010";
ELSIF (OpCode = "10111") THEN	--JC
	q <= "001000011001111100000000010";
ELSIF (OpCode = "11000") THEN	--JMP
	q <= "001000011101111100000000010"; 
ELSIF (OpCode = "11001") THEN	--CALL
	q <= "101000000001000000011100010"; 
ELSIF (OpCode = "11010") THEN	--RET
	q <= "100000000001111100110011001"; 
ELSIF (OpCode = "11011") THEN	--RTI
	q <= "100000000001111100110010101"; 
END IF;
END IF;
END PROCESS;

END a_control_unit;